`timescale 1ps / 1ps
module Filter_Div_31Ux3U_31U_4(
          in2,
          in1,
          out1,
          clk,
          stall
);
   input [30:0] in2;
   input [2:0] in1;
   output [30:0] out1;
   input clk;
   input stall;
wire sub_145_2_n_1, sub_145_2_n_2, sub_145_2_n_3, sub_166_2_n_0, sub_166_2_n_1,
     sub_166_2_n_2, sub_166_2_n_4, sub_187_2_n_0, sub_187_2_n_1, sub_187_2_n_2,
     sub_187_2_n_3, sub_187_2_n_5, sub_187_2_n_7, sub_208_2_n_0, sub_208_2_n_1,
     sub_208_2_n_2, sub_208_2_n_3, sub_208_2_n_5, sub_208_2_n_7, sub_229_2_n_0,
     sub_229_2_n_1, sub_229_2_n_2, sub_229_2_n_3, sub_229_2_n_5, sub_229_2_n_7,
     sub_250_2_n_0, sub_250_2_n_1, sub_250_2_n_2, sub_250_2_n_3, sub_250_2_n_5,
     sub_250_2_n_7, sub_271_2_n_0, sub_271_2_n_1, sub_271_2_n_2, sub_271_2_n_3,
     sub_271_2_n_5, sub_271_2_n_7, sub_292_2_n_0, sub_292_2_n_1, sub_292_2_n_2,
     sub_292_2_n_3, sub_292_2_n_5, sub_292_2_n_7, sub_313_2_n_0, sub_313_2_n_1,
     sub_313_2_n_2, sub_313_2_n_3, sub_313_2_n_5, sub_313_2_n_7, sub_334_2_n_0,
     sub_334_2_n_1, sub_334_2_n_2, sub_334_2_n_3, sub_334_2_n_5, sub_334_2_n_7,
     sub_355_2_n_0, sub_355_2_n_1, sub_355_2_n_2, sub_355_2_n_3, sub_355_2_n_5,
     sub_355_2_n_7, sub_376_2_n_0, sub_376_2_n_1, sub_376_2_n_2, sub_376_2_n_3,
     sub_376_2_n_5, sub_376_2_n_7, sub_397_2_n_0, sub_397_2_n_1, sub_397_2_n_2,
     sub_397_2_n_3, sub_397_2_n_5, sub_397_2_n_7, sub_418_2_n_0, sub_418_2_n_1,
     sub_418_2_n_2, sub_418_2_n_3, sub_418_2_n_5, sub_418_2_n_7, sub_439_2_n_0,
     sub_439_2_n_1, sub_439_2_n_2, sub_439_2_n_3, sub_439_2_n_5, sub_439_2_n_7,
     sub_460_2_n_0, sub_460_2_n_1, sub_460_2_n_2, sub_460_2_n_3, sub_460_2_n_5,
     sub_460_2_n_7, sub_481_2_n_0, sub_481_2_n_1, sub_481_2_n_2, sub_481_2_n_3,
     sub_481_2_n_5, sub_481_2_n_7, sub_502_2_n_0, sub_502_2_n_1, sub_502_2_n_2,
     sub_502_2_n_3, sub_502_2_n_5, sub_502_2_n_7, sub_523_2_n_0, sub_523_2_n_1,
     sub_523_2_n_2, sub_523_2_n_3, sub_523_2_n_5, sub_523_2_n_7, sub_544_2_n_0,
     sub_544_2_n_1, sub_544_2_n_2, sub_544_2_n_3, sub_544_2_n_5, sub_544_2_n_7,
     sub_565_2_n_0, sub_565_2_n_1, sub_565_2_n_2, sub_565_2_n_3, sub_565_2_n_5,
     sub_565_2_n_7, sub_586_2_n_0, sub_586_2_n_1, sub_586_2_n_2, sub_586_2_n_3,
     sub_586_2_n_5, sub_586_2_n_7, sub_607_2_n_0, sub_607_2_n_1, sub_607_2_n_2,
     sub_607_2_n_3, sub_607_2_n_5, sub_607_2_n_7, sub_628_2_n_0, sub_628_2_n_1,
     sub_628_2_n_2, sub_628_2_n_3, sub_628_2_n_5, sub_628_2_n_7, sub_649_2_n_0,
     sub_649_2_n_1, sub_649_2_n_2, sub_649_2_n_3, sub_649_2_n_5, sub_649_2_n_7,
     sub_670_2_n_0, sub_670_2_n_1, sub_670_2_n_2, sub_670_2_n_3, sub_670_2_n_5,
     sub_670_2_n_7, sub_691_2_n_0, sub_691_2_n_1, sub_691_2_n_2, sub_691_2_n_3,
     sub_691_2_n_5, sub_691_2_n_7, sub_712_2_n_0, sub_712_2_n_1, sub_712_2_n_2,
     sub_712_2_n_3, sub_712_2_n_5, sub_712_2_n_7, sub_733_2_n_0, sub_733_2_n_1,
     sub_733_2_n_2, sub_733_2_n_3, sub_733_2_n_5, sub_733_2_n_7, sub_754_2_n_0,
     sub_754_2_n_1, sub_754_2_n_2, sub_754_2_n_3, sub_754_2_n_5, sub_754_2_n_7,
     sub_773_2_n_1, sub_773_2_n_2, sub_773_2_n_3, sub_773_2_n_4, sub_773_2_n_5,
     sub_773_2_n_6, sub_773_2_n_7, stall, clk, n_51, n_52, n_57, n_59, n_71,
     n_72, n_73, n_78, n_79, n_80, n_82, n_83, n_85, n_86, asc001_0_0_,
     asc001_0_1_, asc001_0_2_, asc001_0_3_, asc001_0_4_, asc001_0_5_,
     asc001_0_6_, asc001_0_7_, asc001_0_8_, asc001_0_9_, asc001_0_10_,
     asc001_0_11_, asc001_0_12_, asc001_0_13_, asc001_0_14_, asc001_0_15_,
     asc001_0_16_, asc001_0_17_, asc001_0_18_, asc001_0_19_, asc001_0_20_,
     asc001_0_21_, asc001_0_22_, asc001_0_23_, asc001_0_24_, asc001_0_25_,
     asc001_0_26_, asc001_0_27_, asc001_0_28_, asc001_0_29_, asc001_0_30_,
     in2_1_0_, in2_1_3_, in2_2_0_, in2_4_0_, in2_4_1_, in2_4_3_, in2_5_0_,
     in2_5_1_, in2_7_0_, in2_7_1_, in2_7_2_, in2_7_3_, in2_8_0_, in2_8_1_,
     in2_8_2_, in2_10_0_, in2_10_1_, in2_10_2_, in2_10_3_, in2_11_0_, in2_11_1_,
     in2_11_2_, in2_13_0_, in2_13_1_, in2_13_2_, in2_13_3_, in2_14_0_, in2_14_1_,
     in2_14_2_, in2_16_0_, in2_16_1_, in2_16_2_, in2_16_3_, in2_17_0_, in2_17_1_,
     in2_17_2_, in2_19_0_, in2_19_1_, in2_19_2_, in2_19_3_, in2_20_0_, in2_20_1_,
     in2_20_2_, in2_22_0_, in2_22_1_, in2_22_2_, in2_22_3_, in2_23_0_, in2_23_1_,
     in2_23_2_, in2_25_0_, in2_25_1_, in2_25_2_, in2_25_3_, in2_26_0_, in2_26_1_,
     in2_26_2_, in2_28_0_, in2_28_1_, in2_28_2_, in2_28_3_, in2_29_0_, in2_29_1_,
     in2_29_2_, in2_31_0_, in2_31_1_, in2_31_2_, in2_31_3_, in2_32_0_, in2_32_1_,
     in2_32_2_, in2_34_0_, in2_34_1_, in2_34_2_, in2_34_3_, in2_35_0_, in2_35_1_,
     in2_35_2_, in2_37_0_, in2_37_1_, in2_37_2_, in2_37_3_, in2_38_0_, in2_38_1_,
     in2_38_2_, in2_40_0_, in2_40_1_, in2_40_2_, in2_40_3_, in2_41_0_, in2_41_1_,
     in2_41_2_, in2_43_0_, in2_43_1_, in2_43_2_, in2_43_3_, in2_44_0_, in2_44_1_,
     in2_44_2_, in2_46_0_, in2_46_1_, in2_46_2_, in2_46_3_, in2_47_0_, in2_47_1_,
     in2_47_2_, in2_49_0_, in2_49_1_, in2_49_2_, in2_49_3_, in2_50_0_, in2_50_1_,
     in2_50_2_, in2_52_0_, in2_52_1_, in2_52_2_, in2_52_3_, in2_53_0_, in2_53_1_,
     in2_53_2_, in2_55_0_, in2_55_1_, in2_55_2_, in2_55_3_, in2_56_0_, in2_56_1_,
     in2_56_2_, in2_58_0_, in2_58_1_, in2_58_2_, in2_58_3_, in2_59_0_, in2_59_1_,
     in2_59_2_, in2_61_0_, in2_61_1_, in2_61_2_, in2_61_3_, in2_62_0_, in2_62_1_,
     in2_62_2_, in2_64_0_, in2_64_1_, in2_64_2_, in2_64_3_, in2_65_0_, in2_65_1_,
     in2_65_2_, in2_67_0_, in2_67_1_, in2_67_2_, in2_67_3_, in2_68_0_, in2_68_1_,
     in2_68_2_, in2_70_0_, in2_70_1_, in2_70_2_, in2_70_3_, in2_71_0_, in2_71_1_,
     in2_71_2_, in2_73_0_, in2_73_1_, in2_73_2_, in2_73_3_, in2_74_0_, in2_74_1_,
     in2_74_2_, in2_76_0_, in2_76_1_, in2_76_2_, in2_76_3_, in2_77_0_, in2_77_1_,
     in2_77_2_, in2_79_0_, in2_79_1_, in2_79_2_, in2_79_3_, in2_80_0_, in2_80_1_,
     in2_80_2_, in2_82_0_, in2_82_1_, in2_82_2_, in2_82_3_, in2_83_0_, in2_83_1_,
     in2_83_2_, in2_85_0_, in2_85_1_, in2_85_2_, in2_85_3_, in2_86_0_, in2_86_1_,
     in2_86_2_, in2_88_0_, in2_88_1_, in2_88_2_, in2_88_3_, in2_89_0_, in2_89_1_,
     in2_89_2_, in2_91_3_;
assign {out1[7]} = asc001_0_7_;
assign {out1[6]} = asc001_0_6_;
assign {out1[5]} = asc001_0_5_;
assign {out1[4]} = asc001_0_4_;
assign {out1[3]} = asc001_0_3_;
assign {out1[2]} = asc001_0_2_;
assign {out1[1]} = asc001_0_1_;
assign {out1[0]} = asc001_0_0_;
reg cadence_register_n_51;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_51 <= in1[2];
    end
 end
 assign n_51 = cadence_register_n_51;
reg cadence_register_n_52;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_52 <= in2_68_2_;
    end
 end
 assign n_52 = cadence_register_n_52;
reg cadence_register_out1_8;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_8 <= asc001_0_8_;
    end
 end
 assign out1[8] = cadence_register_out1_8;
reg cadence_register_out1_25;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_25 <= asc001_0_25_;
    end
 end
 assign out1[25] = cadence_register_out1_25;
reg cadence_register_out1_30;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_30 <= asc001_0_30_;
    end
 end
 assign out1[30] = cadence_register_out1_30;
reg cadence_register_out1_23;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_23 <= asc001_0_23_;
    end
 end
 assign out1[23] = cadence_register_out1_23;
reg cadence_register_n_57;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_57 <= in1[0];
    end
 end
 assign n_57 = cadence_register_n_57;
reg cadence_register_out1_10;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_10 <= asc001_0_10_;
    end
 end
 assign out1[10] = cadence_register_out1_10;
reg cadence_register_n_59;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_59 <= sub_773_2_n_5;
    end
 end
 assign n_59 = cadence_register_n_59;
reg cadence_register_out1_11;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_11 <= asc001_0_11_;
    end
 end
 assign out1[11] = cadence_register_out1_11;
reg cadence_register_out1_14;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_14 <= asc001_0_14_;
    end
 end
 assign out1[14] = cadence_register_out1_14;
reg cadence_register_out1_13;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_13 <= asc001_0_13_;
    end
 end
 assign out1[13] = cadence_register_out1_13;
reg cadence_register_out1_12;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_12 <= asc001_0_12_;
    end
 end
 assign out1[12] = cadence_register_out1_12;
reg cadence_register_out1_16;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_16 <= asc001_0_16_;
    end
 end
 assign out1[16] = cadence_register_out1_16;
reg cadence_register_out1_17;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_17 <= asc001_0_17_;
    end
 end
 assign out1[17] = cadence_register_out1_17;
reg cadence_register_out1_20;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_20 <= asc001_0_20_;
    end
 end
 assign out1[20] = cadence_register_out1_20;
reg cadence_register_out1_19;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_19 <= asc001_0_19_;
    end
 end
 assign out1[19] = cadence_register_out1_19;
reg cadence_register_out1_21;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_21 <= asc001_0_21_;
    end
 end
 assign out1[21] = cadence_register_out1_21;
reg cadence_register_out1_22;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_22 <= asc001_0_22_;
    end
 end
 assign out1[22] = cadence_register_out1_22;
reg cadence_register_out1_26;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_26 <= asc001_0_26_;
    end
 end
 assign out1[26] = cadence_register_out1_26;
reg cadence_register_n_71;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_71 <= in1[1];
    end
 end
 assign n_71 = cadence_register_n_71;
reg cadence_register_n_72;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_72 <= in2[2];
    end
 end
 assign n_72 = cadence_register_n_72;
reg cadence_register_n_73;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_73 <= in2_68_0_;
    end
 end
 assign n_73 = cadence_register_n_73;
reg cadence_register_out1_27;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_27 <= asc001_0_27_;
    end
 end
 assign out1[27] = cadence_register_out1_27;
reg cadence_register_out1_24;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_24 <= asc001_0_24_;
    end
 end
 assign out1[24] = cadence_register_out1_24;
reg cadence_register_out1_15;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_15 <= asc001_0_15_;
    end
 end
 assign out1[15] = cadence_register_out1_15;
reg cadence_register_out1_28;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_28 <= asc001_0_28_;
    end
 end
 assign out1[28] = cadence_register_out1_28;
reg cadence_register_n_78;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_78 <= in2[4];
    end
 end
 assign n_78 = cadence_register_n_78;
reg cadence_register_n_79;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_79 <= in2[7];
    end
 end
 assign n_79 = cadence_register_n_79;
reg cadence_register_n_80;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_80 <= in2[6];
    end
 end
 assign n_80 = cadence_register_n_80;
reg cadence_register_out1_29;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_29 <= asc001_0_29_;
    end
 end
 assign out1[29] = cadence_register_out1_29;
reg cadence_register_n_82;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_82 <= in2[5];
    end
 end
 assign n_82 = cadence_register_n_82;
reg cadence_register_n_83;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_83 <= in2_68_1_;
    end
 end
 assign n_83 = cadence_register_n_83;
reg cadence_register_out1_9;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_9 <= asc001_0_9_;
    end
 end
 assign out1[9] = cadence_register_out1_9;
reg cadence_register_n_85;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_85 <= in2[1];
    end
 end
 assign n_85 = cadence_register_n_85;
reg cadence_register_n_86;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_86 <= in2[3];
    end
 end
 assign n_86 = cadence_register_n_86;
reg cadence_register_out1_18;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_18 <= asc001_0_18_;
    end
 end
 assign out1[18] = cadence_register_out1_18;
 assign asc001_0_0_ = ~in2_91_3_;
 assign in2_2_0_ = ((in2_1_0_ & ~in2_1_3_) | ({in2[30]} & in2_1_3_));
 assign in2_5_1_ = ((in2_4_1_ & ~in2_4_3_) | (in2_2_0_ & in2_4_3_));
 assign in2_5_0_ = ((in2_4_0_ & ~in2_4_3_) | ({in2[29]} & in2_4_3_));
 assign in2_8_2_ = ((in2_7_2_ & ~in2_7_3_) | (in2_5_1_ & in2_7_3_));
 assign in2_8_1_ = ((in2_7_1_ & ~in2_7_3_) | (in2_5_0_ & in2_7_3_));
 assign in2_8_0_ = ((in2_7_0_ & ~in2_7_3_) | ({in2[28]} & in2_7_3_));
 assign in2_11_2_ = ((in2_10_2_ & ~in2_10_3_) | (in2_8_1_ & in2_10_3_));
 assign in2_11_1_ = ((in2_10_1_ & ~in2_10_3_) | (in2_8_0_ & in2_10_3_));
 assign in2_11_0_ = ((in2_10_0_ & ~in2_10_3_) | ({in2[27]} & in2_10_3_));
 assign in2_14_2_ = ((in2_13_2_ & ~in2_13_3_) | (in2_11_1_ & in2_13_3_));
 assign in2_14_1_ = ((in2_13_1_ & ~in2_13_3_) | (in2_11_0_ & in2_13_3_));
 assign in2_14_0_ = ((in2_13_0_ & ~in2_13_3_) | ({in2[26]} & in2_13_3_));
 assign in2_17_2_ = ((in2_16_2_ & ~in2_16_3_) | (in2_14_1_ & in2_16_3_));
 assign in2_17_1_ = ((in2_16_1_ & ~in2_16_3_) | (in2_14_0_ & in2_16_3_));
 assign in2_17_0_ = ((in2_16_0_ & ~in2_16_3_) | ({in2[25]} & in2_16_3_));
 assign in2_20_2_ = ((in2_19_2_ & ~in2_19_3_) | (in2_17_1_ & in2_19_3_));
 assign in2_20_1_ = ((in2_19_1_ & ~in2_19_3_) | (in2_17_0_ & in2_19_3_));
 assign in2_20_0_ = ((in2_19_0_ & ~in2_19_3_) | ({in2[24]} & in2_19_3_));
 assign in2_23_2_ = ((in2_22_2_ & ~in2_22_3_) | (in2_20_1_ & in2_22_3_));
 assign in2_23_1_ = ((in2_22_1_ & ~in2_22_3_) | (in2_20_0_ & in2_22_3_));
 assign in2_23_0_ = ((in2_22_0_ & ~in2_22_3_) | ({in2[23]} & in2_22_3_));
 assign in2_26_2_ = ((in2_25_2_ & ~in2_25_3_) | (in2_23_1_ & in2_25_3_));
 assign in2_26_1_ = ((in2_25_1_ & ~in2_25_3_) | (in2_23_0_ & in2_25_3_));
 assign in2_26_0_ = ((in2_25_0_ & ~in2_25_3_) | ({in2[22]} & in2_25_3_));
 assign in2_29_2_ = ((in2_28_2_ & ~in2_28_3_) | (in2_26_1_ & in2_28_3_));
 assign in2_29_1_ = ((in2_28_1_ & ~in2_28_3_) | (in2_26_0_ & in2_28_3_));
 assign in2_29_0_ = ((in2_28_0_ & ~in2_28_3_) | ({in2[21]} & in2_28_3_));
 assign in2_32_2_ = ((in2_31_2_ & ~in2_31_3_) | (in2_29_1_ & in2_31_3_));
 assign in2_32_1_ = ((in2_31_1_ & ~in2_31_3_) | (in2_29_0_ & in2_31_3_));
 assign in2_32_0_ = ((in2_31_0_ & ~in2_31_3_) | ({in2[20]} & in2_31_3_));
 assign in2_35_2_ = ((in2_34_2_ & ~in2_34_3_) | (in2_32_1_ & in2_34_3_));
 assign in2_35_1_ = ((in2_34_1_ & ~in2_34_3_) | (in2_32_0_ & in2_34_3_));
 assign in2_35_0_ = ((in2_34_0_ & ~in2_34_3_) | ({in2[19]} & in2_34_3_));
 assign in2_38_2_ = ((in2_37_2_ & ~in2_37_3_) | (in2_35_1_ & in2_37_3_));
 assign in2_38_1_ = ((in2_37_1_ & ~in2_37_3_) | (in2_35_0_ & in2_37_3_));
 assign in2_38_0_ = ((in2_37_0_ & ~in2_37_3_) | ({in2[18]} & in2_37_3_));
 assign in2_41_2_ = ((in2_40_2_ & ~in2_40_3_) | (in2_38_1_ & in2_40_3_));
 assign in2_41_1_ = ((in2_40_1_ & ~in2_40_3_) | (in2_38_0_ & in2_40_3_));
 assign in2_41_0_ = ((in2_40_0_ & ~in2_40_3_) | ({in2[17]} & in2_40_3_));
 assign in2_44_2_ = ((in2_43_2_ & ~in2_43_3_) | (in2_41_1_ & in2_43_3_));
 assign in2_44_1_ = ((in2_43_1_ & ~in2_43_3_) | (in2_41_0_ & in2_43_3_));
 assign in2_44_0_ = ((in2_43_0_ & ~in2_43_3_) | ({in2[16]} & in2_43_3_));
 assign in2_47_2_ = ((in2_46_2_ & ~in2_46_3_) | (in2_44_1_ & in2_46_3_));
 assign in2_47_1_ = ((in2_46_1_ & ~in2_46_3_) | (in2_44_0_ & in2_46_3_));
 assign in2_47_0_ = ((in2_46_0_ & ~in2_46_3_) | ({in2[15]} & in2_46_3_));
 assign in2_50_2_ = ((in2_49_2_ & ~in2_49_3_) | (in2_47_1_ & in2_49_3_));
 assign in2_50_1_ = ((in2_49_1_ & ~in2_49_3_) | (in2_47_0_ & in2_49_3_));
 assign in2_50_0_ = ((in2_49_0_ & ~in2_49_3_) | ({in2[14]} & in2_49_3_));
 assign in2_53_2_ = ((in2_52_2_ & ~in2_52_3_) | (in2_50_1_ & in2_52_3_));
 assign in2_53_1_ = ((in2_52_1_ & ~in2_52_3_) | (in2_50_0_ & in2_52_3_));
 assign in2_53_0_ = ((in2_52_0_ & ~in2_52_3_) | ({in2[13]} & in2_52_3_));
 assign in2_56_2_ = ((in2_55_2_ & ~in2_55_3_) | (in2_53_1_ & in2_55_3_));
 assign in2_56_1_ = ((in2_55_1_ & ~in2_55_3_) | (in2_53_0_ & in2_55_3_));
 assign in2_56_0_ = ((in2_55_0_ & ~in2_55_3_) | ({in2[12]} & in2_55_3_));
 assign in2_59_2_ = ((in2_58_2_ & ~in2_58_3_) | (in2_56_1_ & in2_58_3_));
 assign in2_59_1_ = ((in2_58_1_ & ~in2_58_3_) | (in2_56_0_ & in2_58_3_));
 assign in2_59_0_ = ((in2_58_0_ & ~in2_58_3_) | ({in2[11]} & in2_58_3_));
 assign in2_62_2_ = ((in2_61_2_ & ~in2_61_3_) | (in2_59_1_ & in2_61_3_));
 assign in2_62_1_ = ((in2_61_1_ & ~in2_61_3_) | (in2_59_0_ & in2_61_3_));
 assign in2_62_0_ = ((in2_61_0_ & ~in2_61_3_) | ({in2[10]} & in2_61_3_));
 assign in2_65_2_ = ((in2_64_2_ & ~in2_64_3_) | (in2_62_1_ & in2_64_3_));
 assign in2_65_1_ = ((in2_64_1_ & ~in2_64_3_) | (in2_62_0_ & in2_64_3_));
 assign in2_65_0_ = ((in2_64_0_ & ~in2_64_3_) | ({in2[9]} & in2_64_3_));
 assign in2_68_2_ = ((in2_67_2_ & ~in2_67_3_) | (in2_65_1_ & in2_67_3_));
 assign in2_68_1_ = ((in2_67_1_ & ~in2_67_3_) | (in2_65_0_ & in2_67_3_));
 assign in2_68_0_ = ((in2_67_0_ & ~in2_67_3_) | ({in2[8]} & in2_67_3_));
 assign in2_71_2_ = ((in2_70_2_ & ~in2_70_3_) | (n_83 & in2_70_3_));
 assign in2_71_1_ = ((in2_70_1_ & ~in2_70_3_) | (n_73 & in2_70_3_));
 assign in2_71_0_ = ((in2_70_0_ & ~in2_70_3_) | (n_79 & in2_70_3_));
 assign in2_74_2_ = ((in2_73_2_ & ~in2_73_3_) | (in2_71_1_ & in2_73_3_));
 assign in2_74_1_ = ((in2_73_1_ & ~in2_73_3_) | (in2_71_0_ & in2_73_3_));
 assign in2_74_0_ = ((in2_73_0_ & ~in2_73_3_) | (n_80 & in2_73_3_));
 assign in2_77_2_ = ((in2_76_2_ & ~in2_76_3_) | (in2_74_1_ & in2_76_3_));
 assign in2_77_1_ = ((in2_76_1_ & ~in2_76_3_) | (in2_74_0_ & in2_76_3_));
 assign in2_77_0_ = ((in2_76_0_ & ~in2_76_3_) | (n_82 & in2_76_3_));
 assign in2_80_2_ = ((in2_79_2_ & ~in2_79_3_) | (in2_77_1_ & in2_79_3_));
 assign in2_80_1_ = ((in2_79_1_ & ~in2_79_3_) | (in2_77_0_ & in2_79_3_));
 assign in2_80_0_ = ((in2_79_0_ & ~in2_79_3_) | (n_78 & in2_79_3_));
 assign in2_83_2_ = ((in2_82_2_ & ~in2_82_3_) | (in2_80_1_ & in2_82_3_));
 assign in2_83_1_ = ((in2_82_1_ & ~in2_82_3_) | (in2_80_0_ & in2_82_3_));
 assign in2_83_0_ = ((in2_82_0_ & ~in2_82_3_) | (n_86 & in2_82_3_));
 assign in2_86_2_ = ((in2_85_2_ & ~in2_85_3_) | (in2_83_1_ & in2_85_3_));
 assign in2_86_1_ = ((in2_85_1_ & ~in2_85_3_) | (in2_83_0_ & in2_85_3_));
 assign in2_86_0_ = ((in2_85_0_ & ~in2_85_3_) | (n_72 & in2_85_3_));
 assign in2_89_2_ = ((in2_88_2_ & ~in2_88_3_) | (in2_86_1_ & in2_88_3_));
 assign in2_89_1_ = ((in2_88_1_ & ~in2_88_3_) | (in2_86_0_ & in2_88_3_));
 assign in2_89_0_ = ((in2_88_0_ & ~in2_88_3_) | (n_85 & in2_88_3_));
 assign asc001_0_6_ = ~in2_73_3_;
 assign asc001_0_1_ = ~in2_88_3_;
 assign asc001_0_2_ = ~in2_85_3_;
 assign asc001_0_3_ = ~in2_82_3_;
 assign asc001_0_4_ = ~in2_79_3_;
 assign asc001_0_5_ = ~in2_76_3_;
 assign asc001_0_30_ = ~in2_1_3_;
 assign asc001_0_7_ = ~in2_70_3_;
 assign asc001_0_8_ = ~in2_67_3_;
 assign asc001_0_9_ = ~in2_64_3_;
 assign asc001_0_10_ = ~in2_61_3_;
 assign asc001_0_11_ = ~in2_58_3_;
 assign asc001_0_12_ = ~in2_55_3_;
 assign asc001_0_13_ = ~in2_52_3_;
 assign asc001_0_29_ = ~in2_4_3_;
 assign asc001_0_15_ = ~in2_46_3_;
 assign asc001_0_16_ = ~in2_43_3_;
 assign asc001_0_17_ = ~in2_40_3_;
 assign asc001_0_18_ = ~in2_37_3_;
 assign asc001_0_19_ = ~in2_34_3_;
 assign asc001_0_20_ = ~in2_31_3_;
 assign asc001_0_21_ = ~in2_28_3_;
 assign asc001_0_22_ = ~in2_25_3_;
 assign asc001_0_23_ = ~in2_22_3_;
 assign asc001_0_24_ = ~in2_19_3_;
 assign asc001_0_25_ = ~in2_16_3_;
 assign asc001_0_26_ = ~in2_13_3_;
 assign asc001_0_27_ = ~in2_10_3_;
 assign asc001_0_28_ = ~in2_7_3_;
 assign asc001_0_14_ = ~in2_49_3_;
 assign in2_1_3_ = (sub_145_2_n_2 | ({in1[1]} | {in1[2]}));
 assign in2_1_0_ = ~sub_145_2_n_3;
 assign sub_145_2_n_2 = (sub_145_2_n_1 & {in1[0]});
 assign sub_145_2_n_3 = (sub_145_2_n_1 ^ {in1[0]});
 assign sub_145_2_n_1 = ~{in2[30]};
 assign in2_4_3_ = ~(sub_166_2_n_4 & ~{in1[2]});
 assign sub_166_2_n_4 = ((sub_166_2_n_2 & in2_2_0_) | ((in2_2_0_ & sub_166_2_n_1) | (sub_166_2_n_1 &
    sub_166_2_n_2)));
 assign in2_4_1_ = (in2_2_0_ ^ (sub_166_2_n_1 ^ sub_166_2_n_2));
 assign in2_4_0_ = ~(sub_166_2_n_2 & ~(sub_166_2_n_0 & {in2[29]}));
 assign sub_166_2_n_2 = ~({in1[0]} & ~{in2[29]});
 assign sub_166_2_n_1 = ~{in1[1]};
 assign sub_166_2_n_0 = ~{in1[0]};
 assign in2_7_3_ = ~sub_187_2_n_7;
 assign sub_187_2_n_7 = ((sub_187_2_n_5 & sub_187_2_n_0) | ((sub_187_2_n_0 & in2_5_1_) | (in2_5_1_ &
    sub_187_2_n_5)));
 assign in2_7_2_ = (sub_187_2_n_0 ^ (in2_5_1_ ^ sub_187_2_n_5));
 assign sub_187_2_n_5 = ((sub_187_2_n_3 & in2_5_0_) | ((in2_5_0_ & sub_187_2_n_2) | (sub_187_2_n_2 &
    sub_187_2_n_3)));
 assign in2_7_1_ = (in2_5_0_ ^ (sub_187_2_n_2 ^ sub_187_2_n_3));
 assign in2_7_0_ = ~(sub_187_2_n_3 & ~(sub_187_2_n_1 & {in2[28]}));
 assign sub_187_2_n_3 = ~({in1[0]} & ~{in2[28]});
 assign sub_187_2_n_2 = ~{in1[1]};
 assign sub_187_2_n_1 = ~{in1[0]};
 assign sub_187_2_n_0 = ~{in1[2]};
 assign in2_10_3_ = ~(sub_208_2_n_7 ^ in2_8_2_);
 assign sub_208_2_n_7 = ((sub_208_2_n_5 & sub_208_2_n_0) | ((sub_208_2_n_0 & in2_8_1_) | (in2_8_1_ &
    sub_208_2_n_5)));
 assign in2_10_2_ = (sub_208_2_n_0 ^ (in2_8_1_ ^ sub_208_2_n_5));
 assign sub_208_2_n_5 = ((sub_208_2_n_3 & in2_8_0_) | ((in2_8_0_ & sub_208_2_n_1) | (sub_208_2_n_1 &
    sub_208_2_n_3)));
 assign in2_10_1_ = (in2_8_0_ ^ (sub_208_2_n_1 ^ sub_208_2_n_3));
 assign in2_10_0_ = ~(sub_208_2_n_3 & ~(sub_208_2_n_2 & {in2[27]}));
 assign sub_208_2_n_3 = ~({in1[0]} & ~{in2[27]});
 assign sub_208_2_n_2 = ~{in1[0]};
 assign sub_208_2_n_1 = ~{in1[1]};
 assign sub_208_2_n_0 = ~{in1[2]};
 assign in2_13_3_ = ~(sub_229_2_n_7 ^ in2_11_2_);
 assign sub_229_2_n_7 = ((sub_229_2_n_5 & sub_229_2_n_0) | ((sub_229_2_n_0 & in2_11_1_) | (in2_11_1_
    & sub_229_2_n_5)));
 assign in2_13_2_ = (sub_229_2_n_0 ^ (in2_11_1_ ^ sub_229_2_n_5));
 assign sub_229_2_n_5 = ((sub_229_2_n_3 & in2_11_0_) | ((in2_11_0_ & sub_229_2_n_1) | (sub_229_2_n_1
    & sub_229_2_n_3)));
 assign in2_13_1_ = (in2_11_0_ ^ (sub_229_2_n_1 ^ sub_229_2_n_3));
 assign in2_13_0_ = ~(sub_229_2_n_3 & ~(sub_229_2_n_2 & {in2[26]}));
 assign sub_229_2_n_3 = ~({in1[0]} & ~{in2[26]});
 assign sub_229_2_n_2 = ~{in1[0]};
 assign sub_229_2_n_1 = ~{in1[1]};
 assign sub_229_2_n_0 = ~{in1[2]};
 assign in2_16_3_ = ~(sub_250_2_n_7 ^ in2_14_2_);
 assign sub_250_2_n_7 = ((sub_250_2_n_5 & sub_250_2_n_0) | ((sub_250_2_n_0 & in2_14_1_) | (in2_14_1_
    & sub_250_2_n_5)));
 assign in2_16_2_ = (sub_250_2_n_0 ^ (in2_14_1_ ^ sub_250_2_n_5));
 assign sub_250_2_n_5 = ((sub_250_2_n_3 & in2_14_0_) | ((in2_14_0_ & sub_250_2_n_1) | (sub_250_2_n_1
    & sub_250_2_n_3)));
 assign in2_16_1_ = (in2_14_0_ ^ (sub_250_2_n_1 ^ sub_250_2_n_3));
 assign in2_16_0_ = ~(sub_250_2_n_3 & ~(sub_250_2_n_2 & {in2[25]}));
 assign sub_250_2_n_3 = ~({in1[0]} & ~{in2[25]});
 assign sub_250_2_n_2 = ~{in1[0]};
 assign sub_250_2_n_1 = ~{in1[1]};
 assign sub_250_2_n_0 = ~{in1[2]};
 assign in2_19_3_ = ~(sub_271_2_n_7 ^ in2_17_2_);
 assign sub_271_2_n_7 = ((sub_271_2_n_5 & sub_271_2_n_0) | ((sub_271_2_n_0 & in2_17_1_) | (in2_17_1_
    & sub_271_2_n_5)));
 assign in2_19_2_ = (sub_271_2_n_0 ^ (in2_17_1_ ^ sub_271_2_n_5));
 assign sub_271_2_n_5 = ((sub_271_2_n_3 & in2_17_0_) | ((in2_17_0_ & sub_271_2_n_1) | (sub_271_2_n_1
    & sub_271_2_n_3)));
 assign in2_19_1_ = (in2_17_0_ ^ (sub_271_2_n_1 ^ sub_271_2_n_3));
 assign in2_19_0_ = ~(sub_271_2_n_3 & ~(sub_271_2_n_2 & {in2[24]}));
 assign sub_271_2_n_3 = ~({in1[0]} & ~{in2[24]});
 assign sub_271_2_n_2 = ~{in1[0]};
 assign sub_271_2_n_1 = ~{in1[1]};
 assign sub_271_2_n_0 = ~{in1[2]};
 assign in2_22_3_ = ~(sub_292_2_n_7 ^ in2_20_2_);
 assign sub_292_2_n_7 = ((sub_292_2_n_5 & sub_292_2_n_0) | ((sub_292_2_n_0 & in2_20_1_) | (in2_20_1_
    & sub_292_2_n_5)));
 assign in2_22_2_ = (sub_292_2_n_0 ^ (in2_20_1_ ^ sub_292_2_n_5));
 assign sub_292_2_n_5 = ((sub_292_2_n_3 & in2_20_0_) | ((in2_20_0_ & sub_292_2_n_1) | (sub_292_2_n_1
    & sub_292_2_n_3)));
 assign in2_22_1_ = (in2_20_0_ ^ (sub_292_2_n_1 ^ sub_292_2_n_3));
 assign in2_22_0_ = ~(sub_292_2_n_3 & ~(sub_292_2_n_2 & {in2[23]}));
 assign sub_292_2_n_3 = ~({in1[0]} & ~{in2[23]});
 assign sub_292_2_n_2 = ~{in1[0]};
 assign sub_292_2_n_1 = ~{in1[1]};
 assign sub_292_2_n_0 = ~{in1[2]};
 assign in2_25_3_ = ~(sub_313_2_n_7 ^ in2_23_2_);
 assign sub_313_2_n_7 = ((sub_313_2_n_5 & sub_313_2_n_0) | ((sub_313_2_n_0 & in2_23_1_) | (in2_23_1_
    & sub_313_2_n_5)));
 assign in2_25_2_ = (sub_313_2_n_0 ^ (in2_23_1_ ^ sub_313_2_n_5));
 assign sub_313_2_n_5 = ((sub_313_2_n_3 & in2_23_0_) | ((in2_23_0_ & sub_313_2_n_1) | (sub_313_2_n_1
    & sub_313_2_n_3)));
 assign in2_25_1_ = (in2_23_0_ ^ (sub_313_2_n_1 ^ sub_313_2_n_3));
 assign in2_25_0_ = ~(sub_313_2_n_3 & ~(sub_313_2_n_2 & {in2[22]}));
 assign sub_313_2_n_3 = ~({in1[0]} & ~{in2[22]});
 assign sub_313_2_n_2 = ~{in1[0]};
 assign sub_313_2_n_1 = ~{in1[1]};
 assign sub_313_2_n_0 = ~{in1[2]};
 assign in2_28_3_ = ~(sub_334_2_n_7 ^ in2_26_2_);
 assign sub_334_2_n_7 = ((sub_334_2_n_5 & sub_334_2_n_0) | ((sub_334_2_n_0 & in2_26_1_) | (in2_26_1_
    & sub_334_2_n_5)));
 assign in2_28_2_ = (sub_334_2_n_0 ^ (in2_26_1_ ^ sub_334_2_n_5));
 assign sub_334_2_n_5 = ((sub_334_2_n_3 & in2_26_0_) | ((in2_26_0_ & sub_334_2_n_1) | (sub_334_2_n_1
    & sub_334_2_n_3)));
 assign in2_28_1_ = (in2_26_0_ ^ (sub_334_2_n_1 ^ sub_334_2_n_3));
 assign in2_28_0_ = ~(sub_334_2_n_3 & ~(sub_334_2_n_2 & {in2[21]}));
 assign sub_334_2_n_3 = ~({in1[0]} & ~{in2[21]});
 assign sub_334_2_n_2 = ~{in1[0]};
 assign sub_334_2_n_1 = ~{in1[1]};
 assign sub_334_2_n_0 = ~{in1[2]};
 assign in2_31_3_ = ~(sub_355_2_n_7 ^ in2_29_2_);
 assign sub_355_2_n_7 = ((sub_355_2_n_5 & sub_355_2_n_0) | ((sub_355_2_n_0 & in2_29_1_) | (in2_29_1_
    & sub_355_2_n_5)));
 assign in2_31_2_ = (sub_355_2_n_0 ^ (in2_29_1_ ^ sub_355_2_n_5));
 assign sub_355_2_n_5 = ((sub_355_2_n_3 & in2_29_0_) | ((in2_29_0_ & sub_355_2_n_1) | (sub_355_2_n_1
    & sub_355_2_n_3)));
 assign in2_31_1_ = (in2_29_0_ ^ (sub_355_2_n_1 ^ sub_355_2_n_3));
 assign in2_31_0_ = ~(sub_355_2_n_3 & ~(sub_355_2_n_2 & {in2[20]}));
 assign sub_355_2_n_3 = ~({in1[0]} & ~{in2[20]});
 assign sub_355_2_n_2 = ~{in1[0]};
 assign sub_355_2_n_1 = ~{in1[1]};
 assign sub_355_2_n_0 = ~{in1[2]};
 assign in2_34_3_ = ~(sub_376_2_n_7 ^ in2_32_2_);
 assign sub_376_2_n_7 = ((sub_376_2_n_5 & sub_376_2_n_0) | ((sub_376_2_n_0 & in2_32_1_) | (in2_32_1_
    & sub_376_2_n_5)));
 assign in2_34_2_ = (sub_376_2_n_0 ^ (in2_32_1_ ^ sub_376_2_n_5));
 assign sub_376_2_n_5 = ((sub_376_2_n_3 & in2_32_0_) | ((in2_32_0_ & sub_376_2_n_1) | (sub_376_2_n_1
    & sub_376_2_n_3)));
 assign in2_34_1_ = (in2_32_0_ ^ (sub_376_2_n_1 ^ sub_376_2_n_3));
 assign in2_34_0_ = ~(sub_376_2_n_3 & ~(sub_376_2_n_2 & {in2[19]}));
 assign sub_376_2_n_3 = ~({in1[0]} & ~{in2[19]});
 assign sub_376_2_n_2 = ~{in1[0]};
 assign sub_376_2_n_1 = ~{in1[1]};
 assign sub_376_2_n_0 = ~{in1[2]};
 assign in2_37_3_ = ~(sub_397_2_n_7 ^ in2_35_2_);
 assign sub_397_2_n_7 = ((sub_397_2_n_5 & sub_397_2_n_0) | ((sub_397_2_n_0 & in2_35_1_) | (in2_35_1_
    & sub_397_2_n_5)));
 assign in2_37_2_ = (sub_397_2_n_0 ^ (in2_35_1_ ^ sub_397_2_n_5));
 assign sub_397_2_n_5 = ((sub_397_2_n_3 & in2_35_0_) | ((in2_35_0_ & sub_397_2_n_1) | (sub_397_2_n_1
    & sub_397_2_n_3)));
 assign in2_37_1_ = (in2_35_0_ ^ (sub_397_2_n_1 ^ sub_397_2_n_3));
 assign in2_37_0_ = ~(sub_397_2_n_3 & ~(sub_397_2_n_2 & {in2[18]}));
 assign sub_397_2_n_3 = ~({in1[0]} & ~{in2[18]});
 assign sub_397_2_n_2 = ~{in1[0]};
 assign sub_397_2_n_1 = ~{in1[1]};
 assign sub_397_2_n_0 = ~{in1[2]};
 assign in2_40_3_ = ~(sub_418_2_n_7 ^ in2_38_2_);
 assign sub_418_2_n_7 = ((sub_418_2_n_5 & sub_418_2_n_0) | ((sub_418_2_n_0 & in2_38_1_) | (in2_38_1_
    & sub_418_2_n_5)));
 assign in2_40_2_ = (sub_418_2_n_0 ^ (in2_38_1_ ^ sub_418_2_n_5));
 assign sub_418_2_n_5 = ((sub_418_2_n_3 & in2_38_0_) | ((in2_38_0_ & sub_418_2_n_1) | (sub_418_2_n_1
    & sub_418_2_n_3)));
 assign in2_40_1_ = (in2_38_0_ ^ (sub_418_2_n_1 ^ sub_418_2_n_3));
 assign in2_40_0_ = ~(sub_418_2_n_3 & ~(sub_418_2_n_2 & {in2[17]}));
 assign sub_418_2_n_3 = ~({in1[0]} & ~{in2[17]});
 assign sub_418_2_n_2 = ~{in1[0]};
 assign sub_418_2_n_1 = ~{in1[1]};
 assign sub_418_2_n_0 = ~{in1[2]};
 assign in2_43_3_ = ~(sub_439_2_n_7 ^ in2_41_2_);
 assign sub_439_2_n_7 = ((sub_439_2_n_5 & sub_439_2_n_0) | ((sub_439_2_n_0 & in2_41_1_) | (in2_41_1_
    & sub_439_2_n_5)));
 assign in2_43_2_ = (sub_439_2_n_0 ^ (in2_41_1_ ^ sub_439_2_n_5));
 assign sub_439_2_n_5 = ((sub_439_2_n_3 & in2_41_0_) | ((in2_41_0_ & sub_439_2_n_1) | (sub_439_2_n_1
    & sub_439_2_n_3)));
 assign in2_43_1_ = (in2_41_0_ ^ (sub_439_2_n_1 ^ sub_439_2_n_3));
 assign in2_43_0_ = ~(sub_439_2_n_3 & ~(sub_439_2_n_2 & {in2[16]}));
 assign sub_439_2_n_3 = ~({in1[0]} & ~{in2[16]});
 assign sub_439_2_n_2 = ~{in1[0]};
 assign sub_439_2_n_1 = ~{in1[1]};
 assign sub_439_2_n_0 = ~{in1[2]};
 assign in2_46_3_ = ~(sub_460_2_n_7 ^ in2_44_2_);
 assign sub_460_2_n_7 = ((sub_460_2_n_5 & sub_460_2_n_0) | ((sub_460_2_n_0 & in2_44_1_) | (in2_44_1_
    & sub_460_2_n_5)));
 assign in2_46_2_ = (sub_460_2_n_0 ^ (in2_44_1_ ^ sub_460_2_n_5));
 assign sub_460_2_n_5 = ((sub_460_2_n_3 & in2_44_0_) | ((in2_44_0_ & sub_460_2_n_1) | (sub_460_2_n_1
    & sub_460_2_n_3)));
 assign in2_46_1_ = (in2_44_0_ ^ (sub_460_2_n_1 ^ sub_460_2_n_3));
 assign in2_46_0_ = ~(sub_460_2_n_3 & ~(sub_460_2_n_2 & {in2[15]}));
 assign sub_460_2_n_3 = ~({in1[0]} & ~{in2[15]});
 assign sub_460_2_n_2 = ~{in1[0]};
 assign sub_460_2_n_1 = ~{in1[1]};
 assign sub_460_2_n_0 = ~{in1[2]};
 assign in2_49_3_ = ~(sub_481_2_n_7 ^ in2_47_2_);
 assign sub_481_2_n_7 = ((sub_481_2_n_5 & sub_481_2_n_0) | ((sub_481_2_n_0 & in2_47_1_) | (in2_47_1_
    & sub_481_2_n_5)));
 assign in2_49_2_ = (sub_481_2_n_0 ^ (in2_47_1_ ^ sub_481_2_n_5));
 assign sub_481_2_n_5 = ((sub_481_2_n_3 & in2_47_0_) | ((in2_47_0_ & sub_481_2_n_1) | (sub_481_2_n_1
    & sub_481_2_n_3)));
 assign in2_49_1_ = (in2_47_0_ ^ (sub_481_2_n_1 ^ sub_481_2_n_3));
 assign in2_49_0_ = ~(sub_481_2_n_3 & ~(sub_481_2_n_2 & {in2[14]}));
 assign sub_481_2_n_3 = ~({in1[0]} & ~{in2[14]});
 assign sub_481_2_n_2 = ~{in1[0]};
 assign sub_481_2_n_1 = ~{in1[1]};
 assign sub_481_2_n_0 = ~{in1[2]};
 assign in2_52_3_ = ~(sub_502_2_n_7 ^ in2_50_2_);
 assign sub_502_2_n_7 = ((sub_502_2_n_5 & sub_502_2_n_0) | ((sub_502_2_n_0 & in2_50_1_) | (in2_50_1_
    & sub_502_2_n_5)));
 assign in2_52_2_ = (sub_502_2_n_0 ^ (in2_50_1_ ^ sub_502_2_n_5));
 assign sub_502_2_n_5 = ((sub_502_2_n_3 & in2_50_0_) | ((in2_50_0_ & sub_502_2_n_1) | (sub_502_2_n_1
    & sub_502_2_n_3)));
 assign in2_52_1_ = (in2_50_0_ ^ (sub_502_2_n_1 ^ sub_502_2_n_3));
 assign in2_52_0_ = ~(sub_502_2_n_3 & ~(sub_502_2_n_2 & {in2[13]}));
 assign sub_502_2_n_3 = ~({in1[0]} & ~{in2[13]});
 assign sub_502_2_n_2 = ~{in1[0]};
 assign sub_502_2_n_1 = ~{in1[1]};
 assign sub_502_2_n_0 = ~{in1[2]};
 assign in2_55_3_ = ~(sub_523_2_n_7 ^ in2_53_2_);
 assign sub_523_2_n_7 = ((sub_523_2_n_5 & sub_523_2_n_0) | ((sub_523_2_n_0 & in2_53_1_) | (in2_53_1_
    & sub_523_2_n_5)));
 assign in2_55_2_ = (sub_523_2_n_0 ^ (in2_53_1_ ^ sub_523_2_n_5));
 assign sub_523_2_n_5 = ((sub_523_2_n_3 & in2_53_0_) | ((in2_53_0_ & sub_523_2_n_1) | (sub_523_2_n_1
    & sub_523_2_n_3)));
 assign in2_55_1_ = (in2_53_0_ ^ (sub_523_2_n_1 ^ sub_523_2_n_3));
 assign in2_55_0_ = ~(sub_523_2_n_3 & ~(sub_523_2_n_2 & {in2[12]}));
 assign sub_523_2_n_3 = ~({in1[0]} & ~{in2[12]});
 assign sub_523_2_n_2 = ~{in1[0]};
 assign sub_523_2_n_1 = ~{in1[1]};
 assign sub_523_2_n_0 = ~{in1[2]};
 assign in2_58_3_ = ~(sub_544_2_n_7 ^ in2_56_2_);
 assign sub_544_2_n_7 = ((sub_544_2_n_5 & sub_544_2_n_0) | ((sub_544_2_n_0 & in2_56_1_) | (in2_56_1_
    & sub_544_2_n_5)));
 assign in2_58_2_ = (sub_544_2_n_0 ^ (in2_56_1_ ^ sub_544_2_n_5));
 assign sub_544_2_n_5 = ((sub_544_2_n_3 & in2_56_0_) | ((in2_56_0_ & sub_544_2_n_1) | (sub_544_2_n_1
    & sub_544_2_n_3)));
 assign in2_58_1_ = (in2_56_0_ ^ (sub_544_2_n_1 ^ sub_544_2_n_3));
 assign in2_58_0_ = ~(sub_544_2_n_3 & ~(sub_544_2_n_2 & {in2[11]}));
 assign sub_544_2_n_3 = ~({in1[0]} & ~{in2[11]});
 assign sub_544_2_n_2 = ~{in1[0]};
 assign sub_544_2_n_1 = ~{in1[1]};
 assign sub_544_2_n_0 = ~{in1[2]};
 assign in2_61_3_ = ~(sub_565_2_n_7 ^ in2_59_2_);
 assign sub_565_2_n_7 = ((sub_565_2_n_5 & sub_565_2_n_0) | ((sub_565_2_n_0 & in2_59_1_) | (in2_59_1_
    & sub_565_2_n_5)));
 assign in2_61_2_ = (sub_565_2_n_0 ^ (in2_59_1_ ^ sub_565_2_n_5));
 assign sub_565_2_n_5 = ((sub_565_2_n_3 & in2_59_0_) | ((in2_59_0_ & sub_565_2_n_1) | (sub_565_2_n_1
    & sub_565_2_n_3)));
 assign in2_61_1_ = (in2_59_0_ ^ (sub_565_2_n_1 ^ sub_565_2_n_3));
 assign in2_61_0_ = ~(sub_565_2_n_3 & ~(sub_565_2_n_2 & {in2[10]}));
 assign sub_565_2_n_3 = ~({in1[0]} & ~{in2[10]});
 assign sub_565_2_n_2 = ~{in1[0]};
 assign sub_565_2_n_1 = ~{in1[1]};
 assign sub_565_2_n_0 = ~{in1[2]};
 assign in2_64_3_ = ~(sub_586_2_n_7 ^ in2_62_2_);
 assign sub_586_2_n_7 = ((sub_586_2_n_5 & sub_586_2_n_0) | ((sub_586_2_n_0 & in2_62_1_) | (in2_62_1_
    & sub_586_2_n_5)));
 assign in2_64_2_ = (sub_586_2_n_0 ^ (in2_62_1_ ^ sub_586_2_n_5));
 assign sub_586_2_n_5 = ((sub_586_2_n_3 & in2_62_0_) | ((in2_62_0_ & sub_586_2_n_1) | (sub_586_2_n_1
    & sub_586_2_n_3)));
 assign in2_64_1_ = (in2_62_0_ ^ (sub_586_2_n_1 ^ sub_586_2_n_3));
 assign in2_64_0_ = ~(sub_586_2_n_3 & ~(sub_586_2_n_2 & {in2[9]}));
 assign sub_586_2_n_3 = ~({in1[0]} & ~{in2[9]});
 assign sub_586_2_n_2 = ~{in1[0]};
 assign sub_586_2_n_1 = ~{in1[1]};
 assign sub_586_2_n_0 = ~{in1[2]};
 assign in2_67_3_ = ~(sub_607_2_n_7 ^ in2_65_2_);
 assign sub_607_2_n_7 = ((sub_607_2_n_5 & sub_607_2_n_0) | ((sub_607_2_n_0 & in2_65_1_) | (in2_65_1_
    & sub_607_2_n_5)));
 assign in2_67_2_ = (sub_607_2_n_0 ^ (in2_65_1_ ^ sub_607_2_n_5));
 assign sub_607_2_n_5 = ((sub_607_2_n_3 & in2_65_0_) | ((in2_65_0_ & sub_607_2_n_1) | (sub_607_2_n_1
    & sub_607_2_n_3)));
 assign in2_67_1_ = (in2_65_0_ ^ (sub_607_2_n_1 ^ sub_607_2_n_3));
 assign in2_67_0_ = ~(sub_607_2_n_3 & ~(sub_607_2_n_2 & {in2[8]}));
 assign sub_607_2_n_3 = ~({in1[0]} & ~{in2[8]});
 assign sub_607_2_n_2 = ~{in1[0]};
 assign sub_607_2_n_1 = ~{in1[1]};
 assign sub_607_2_n_0 = ~{in1[2]};
 assign in2_70_3_ = ~(sub_628_2_n_7 ^ n_52);
 assign sub_628_2_n_7 = ((sub_628_2_n_5 & sub_628_2_n_0) | ((sub_628_2_n_0 & n_83) | (n_83 & sub_628_2_n_5)));
 assign in2_70_2_ = (sub_628_2_n_0 ^ (n_83 ^ sub_628_2_n_5));
 assign sub_628_2_n_5 = ((sub_628_2_n_3 & n_73) | ((n_73 & sub_628_2_n_1) | (sub_628_2_n_1 & sub_628_2_n_3)));
 assign in2_70_1_ = (n_73 ^ (sub_628_2_n_1 ^ sub_628_2_n_3));
 assign in2_70_0_ = ~(sub_628_2_n_3 & ~(sub_628_2_n_2 & n_79));
 assign sub_628_2_n_3 = ~(n_57 & ~n_79);
 assign sub_628_2_n_2 = ~n_57;
 assign sub_628_2_n_1 = ~n_71;
 assign sub_628_2_n_0 = ~n_51;
 assign in2_73_3_ = ~(sub_649_2_n_7 ^ in2_71_2_);
 assign sub_649_2_n_7 = ((sub_649_2_n_5 & sub_649_2_n_0) | ((sub_649_2_n_0 & in2_71_1_) | (in2_71_1_
    & sub_649_2_n_5)));
 assign in2_73_2_ = (sub_649_2_n_0 ^ (in2_71_1_ ^ sub_649_2_n_5));
 assign sub_649_2_n_5 = ((sub_649_2_n_3 & in2_71_0_) | ((in2_71_0_ & sub_649_2_n_1) | (sub_649_2_n_1
    & sub_649_2_n_3)));
 assign in2_73_1_ = (in2_71_0_ ^ (sub_649_2_n_1 ^ sub_649_2_n_3));
 assign in2_73_0_ = ~(sub_649_2_n_3 & ~(sub_649_2_n_2 & n_80));
 assign sub_649_2_n_3 = ~(n_57 & ~n_80);
 assign sub_649_2_n_2 = ~n_57;
 assign sub_649_2_n_1 = ~n_71;
 assign sub_649_2_n_0 = ~n_51;
 assign in2_76_3_ = ~(sub_670_2_n_7 ^ in2_74_2_);
 assign sub_670_2_n_7 = ((sub_670_2_n_5 & sub_670_2_n_0) | ((sub_670_2_n_0 & in2_74_1_) | (in2_74_1_
    & sub_670_2_n_5)));
 assign in2_76_2_ = (sub_670_2_n_0 ^ (in2_74_1_ ^ sub_670_2_n_5));
 assign sub_670_2_n_5 = ((sub_670_2_n_3 & in2_74_0_) | ((in2_74_0_ & sub_670_2_n_1) | (sub_670_2_n_1
    & sub_670_2_n_3)));
 assign in2_76_1_ = (in2_74_0_ ^ (sub_670_2_n_1 ^ sub_670_2_n_3));
 assign in2_76_0_ = ~(sub_670_2_n_3 & ~(sub_670_2_n_2 & n_82));
 assign sub_670_2_n_3 = ~(n_57 & ~n_82);
 assign sub_670_2_n_2 = ~n_57;
 assign sub_670_2_n_1 = ~n_71;
 assign sub_670_2_n_0 = ~n_51;
 assign in2_79_3_ = ~(sub_691_2_n_7 ^ in2_77_2_);
 assign sub_691_2_n_7 = ((sub_691_2_n_5 & sub_691_2_n_0) | ((sub_691_2_n_0 & in2_77_1_) | (in2_77_1_
    & sub_691_2_n_5)));
 assign in2_79_2_ = (sub_691_2_n_0 ^ (in2_77_1_ ^ sub_691_2_n_5));
 assign sub_691_2_n_5 = ((sub_691_2_n_3 & in2_77_0_) | ((in2_77_0_ & sub_691_2_n_1) | (sub_691_2_n_1
    & sub_691_2_n_3)));
 assign in2_79_1_ = (in2_77_0_ ^ (sub_691_2_n_1 ^ sub_691_2_n_3));
 assign in2_79_0_ = ~(sub_691_2_n_3 & ~(sub_691_2_n_2 & n_78));
 assign sub_691_2_n_3 = ~(n_57 & ~n_78);
 assign sub_691_2_n_2 = ~n_57;
 assign sub_691_2_n_1 = ~n_71;
 assign sub_691_2_n_0 = ~n_51;
 assign in2_82_3_ = ~(sub_712_2_n_7 ^ in2_80_2_);
 assign sub_712_2_n_7 = ((sub_712_2_n_5 & sub_712_2_n_0) | ((sub_712_2_n_0 & in2_80_1_) | (in2_80_1_
    & sub_712_2_n_5)));
 assign in2_82_2_ = (sub_712_2_n_0 ^ (in2_80_1_ ^ sub_712_2_n_5));
 assign sub_712_2_n_5 = ((sub_712_2_n_3 & in2_80_0_) | ((in2_80_0_ & sub_712_2_n_1) | (sub_712_2_n_1
    & sub_712_2_n_3)));
 assign in2_82_1_ = (in2_80_0_ ^ (sub_712_2_n_1 ^ sub_712_2_n_3));
 assign in2_82_0_ = ~(sub_712_2_n_3 & ~(sub_712_2_n_2 & n_86));
 assign sub_712_2_n_3 = ~(n_57 & ~n_86);
 assign sub_712_2_n_2 = ~n_57;
 assign sub_712_2_n_1 = ~n_71;
 assign sub_712_2_n_0 = ~n_51;
 assign in2_85_3_ = ~(sub_733_2_n_7 ^ in2_83_2_);
 assign sub_733_2_n_7 = ((sub_733_2_n_5 & sub_733_2_n_0) | ((sub_733_2_n_0 & in2_83_1_) | (in2_83_1_
    & sub_733_2_n_5)));
 assign in2_85_2_ = (sub_733_2_n_0 ^ (in2_83_1_ ^ sub_733_2_n_5));
 assign sub_733_2_n_5 = ((sub_733_2_n_3 & in2_83_0_) | ((in2_83_0_ & sub_733_2_n_1) | (sub_733_2_n_1
    & sub_733_2_n_3)));
 assign in2_85_1_ = (in2_83_0_ ^ (sub_733_2_n_1 ^ sub_733_2_n_3));
 assign in2_85_0_ = ~(sub_733_2_n_3 & ~(sub_733_2_n_2 & n_72));
 assign sub_733_2_n_3 = ~(n_57 & ~n_72);
 assign sub_733_2_n_2 = ~n_57;
 assign sub_733_2_n_1 = ~n_71;
 assign sub_733_2_n_0 = ~n_51;
 assign in2_88_3_ = ~(sub_754_2_n_7 ^ in2_86_2_);
 assign sub_754_2_n_7 = ((sub_754_2_n_5 & sub_754_2_n_0) | ((sub_754_2_n_0 & in2_86_1_) | (in2_86_1_
    & sub_754_2_n_5)));
 assign in2_88_2_ = (sub_754_2_n_0 ^ (in2_86_1_ ^ sub_754_2_n_5));
 assign sub_754_2_n_5 = ((sub_754_2_n_3 & in2_86_0_) | ((in2_86_0_ & sub_754_2_n_1) | (sub_754_2_n_1
    & sub_754_2_n_3)));
 assign in2_88_1_ = (in2_86_0_ ^ (sub_754_2_n_1 ^ sub_754_2_n_3));
 assign in2_88_0_ = ~(sub_754_2_n_3 & ~(sub_754_2_n_2 & n_85));
 assign sub_754_2_n_3 = ~(n_57 & ~n_85);
 assign sub_754_2_n_2 = ~n_57;
 assign sub_754_2_n_1 = ~n_71;
 assign sub_754_2_n_0 = ~n_51;
 assign in2_91_3_ = ~(sub_773_2_n_7 ^ in2_89_2_);
 assign sub_773_2_n_7 = ~((sub_773_2_n_6 | sub_773_2_n_4) & (n_51 | sub_773_2_n_2));
 assign sub_773_2_n_6 = ~((n_59 & sub_773_2_n_3) | (sub_773_2_n_1 & in2_89_0_));
 assign sub_773_2_n_5 = ~({in1[0]} & ~{in2[0]});
 assign sub_773_2_n_4 = ~(in2_89_1_ | ~n_51);
 assign sub_773_2_n_3 = (in2_89_0_ | sub_773_2_n_1);
 assign sub_773_2_n_2 = ~in2_89_1_;
 assign sub_773_2_n_1 = ~n_71;
endmodule

